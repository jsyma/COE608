library verilog;
use verilog.vl_types.all;
entity lab3_block_vlg_vec_tst is
end lab3_block_vlg_vec_tst;
