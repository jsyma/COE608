library ieee;
use ieee.std_logic_1164.all;

entity bufr is 
port(
	A	:	IN STD_LOGIC_VECTOR(3 downto 0);
	B	:	IN STD_LOGIC_VECTOR(3 downto 0);
	outA	: OUT STD_LOGIC_VECTOR(31 downto 0);
	outB	:	OUT STD_LOGIC_VECTOR(31 downto 0)
);
end bufr;

architecture Behavior of bufr is
begin
	outA <=  "00000000000000000000000000000000" when A = "0000" else
				"00000000000000000000000000000001" when A = "0001" else
				"00000000000000000000000000000010" when A = "0010" else
				"00000000000000000000000000000011" when A = "0011" else
				"00000000000000000000000000000100" when A = "0100" else
				"00000000000000000000000000000101" when A = "0101" else
				"00000000000000000000000000000110" when A = "0110" else
				"00000000000000000000000000000111" when A = "0111" else
				"00000000000000000000000000001000" when A = "1000" else
				"00000000000000000000000000001001" when A = "1001" else
				"00000000000000000000000000001010" when A = "1010" else
				"00000000000000000000000000001011" when A = "1011" else
				"00000000000000000000000000001100" when A = "1100" else
				"00000000000000000000000000001101" when A = "1101" else
				"00000000000000000000000000001110" when A = "1110" else
				"00000000000000000000000000001111" when A = "1111" else
				"00000000000000000000000000000000";
	outB <=  "00000000000000000000000000000000" when B = "0000" else
				"00000000000000000000000000000001" when B = "0001" else
				"00000000000000000000000000000010" when B = "0010" else
				"00000000000000000000000000000011" when B = "0011" else
				"00000000000000000000000000000100" when B = "0100" else
				"00000000000000000000000000000101" when B = "0101" else
				"00000000000000000000000000000110" when B = "0110" else
				"00000000000000000000000000000111" when B = "0111" else
				"00000000000000000000000000001000" when B = "1000" else
				"00000000000000000000000000001001" when B = "1001" else
				"00000000000000000000000000001010" when B = "1010" else
				"00000000000000000000000000001011" when B = "1011" else
				"00000000000000000000000000001100" when B = "1100" else
				"00000000000000000000000000001101" when B = "1101" else
				"00000000000000000000000000001110" when B = "1110" else
				"00000000000000000000000000001111" when B = "1111" else
				"00000000000000000000000000000000";
	
end Behavior;

